
module virtual_IO_16 (
	source,
	probe);	

	output	[15:0]	source;
	input	[15:0]	probe;
endmodule
