// virtualprobe_16bit.v

// Generated using ACDS version 22.1 917

`timescale 1 ps / 1 ps
module virtualprobe_16bit #(NAME="NONE") (
		input  wire [15:0] probe  // probes.probe
	);

	altsource_probe_top #(
		.sld_auto_instance_index ("YES"),
		.sld_instance_index      (0),
		.instance_id             (NAME),
		.probe_width             (16),
		.source_width            (0),
		.enable_metastability    ("NO")
	) in_system_sources_probes_0 (
		.probe (probe)  // probes.probe
	);

endmodule
