
module virtualprobe_16bit (
	probe);	

	input	[15:0]	probe;
endmodule
