//TODO.  need to work out this
module via(clk, rst_n, enable, reg_select, data_bus , porta, portb);
    input clk;
    input rst_n;
    input enable;
    input [3:0] reg_select;
    inout [7:0] data_bus;
    inout [7:0] porta;
    inout [7:0] portb;



endmodule